* C:\Users\admin\Desktop\FOSSEE\parity_checker.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/15/21 21:26:06

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ parity_checker		
U2  Net-_R1-Pad2_ Net-_U1-Pad1_ adc_bridge_1		
U3  Net-_U1-Pad2_ Net-_R2-Pad2_ dac_bridge_1		
R1  Net-_R1-Pad1_ Net-_R1-Pad2_ 100k		
R2  Net-_R1-Pad1_ Net-_R2-Pad2_ 100k		
v1  Net-_R1-Pad2_ Net-_R1-Pad1_ pulse		

.end
